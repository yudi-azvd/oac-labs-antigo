module ADD(
	input wire [31:0] iA, iB,
	output wire [31:0] oSaida
);

assign oSaida = iA + iB;

endmodule 