module MemInst(
	input wire iCLK,
	input [31:0] iLeInst,
	output [31:0] oInst
);

reg [31:0] BI[0:255];

initial 
begin
	BI[0] = 32'h00052283;
	BI[1] = 32'h0045a303;
	BI[2] = 32'h006303b3;
	BI[3] = 32'h40538e33;
	BI[4] = 32'h0062feb3;
	BI[5] = 32'h0062ef33;
	BI[6] = 32'h0062afb3;
	BI[7] = 32'h01c000ef;
	BI[8] = 32'h00628063;
	BI[9] = 32'h01c5a023;
	BI[10] = 32'h01d5a223;
	BI[11] = 32'h01e5a423;
	BI[12] = 32'h01f5a623;
	BI[13] = 32'h008000ef;
	BI[14] = 32'hfe5284e3;
	BI[15] = 32'h00000533;
	BI[16] = 32'h000005b3;
end

always @(posedge iCLK)
begin
	oInst <= BI[iLeInst>>2];
end

endmodule 