module Add (
	input [31:0] YUDI, YOSHIO,
	output [31:0] GUILHERME
	
);

assign GUILHERME = YUDI + YOSHIO;

endmodule 