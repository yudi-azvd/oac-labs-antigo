module AND (
	input iA, iB,
	output oSaida
);

	assign oSaida = iA & iB;

endmodule 